/**
* alu: ALU result
* mem: Data read from the data memory
*/
module cpu (clock, resetn, inst, mem, pc, wmem, alu, data);
   input [31:0] inst, mem;
   input clock, resetn;
   output [31:0] pc, alu, data;
   output wmem;

   wire [31:0]   p4, bpc,
      npc,     // Next value of the PC, selected from 4 inputs
      adr,
      ra,      // 1st value read from the register file
      alua, alub,
      res,     // Data to write to the register
      // ALU result or the data read from the data memory
      alu_mem;
   wire [3:0]    aluc;                 // ALU control signals

   // The number of the register to be written to, either rt or rd
   wire [4:0]    reg_dest,
      // The number of the register to be written to, selected from reg_dest
      // and $ra
      wn;   
   wire [1:0]    pcsource;
   
   // signals generated by CU
   wire wmem, wreg, regrt, m2reg, shift, aluimm, jal, sext;
   wire zero;  // zero flag of ALU

   // extend the immediate value
   wire          e = sext & inst[15];          // positive or negative sign at sext signal
   wire [15:0]   imm = {16{e}};                // high 16 sign bit
   wire [31:0]   immediate = {imm, inst[15:0]};    // sign-extended immediate value

   // shift amount, extended to 32 bits
   wire [31:0]   sa = { 27'b0, inst[10:6] };
   // branch offset
   wire [31:0]   offset = {imm[13:0], inst[15:0], 1'b0, 1'b0};

   dff32 ip (npc, clock, resetn, pc);  // define a D-register for PC
   
   // cla32 pcplus4 (pc, 32'h4, 1'b0, p4);
   // cla32 br_adr (p4, offset, 1'b0, adr);
   
   assign p4 = pc + 32'h4;       // modified
   assign adr = p4 + offset;     // branch address
   
   wire [31:0] jpc = {p4[31:28], inst[25:0], 2'b00}; // j address 
   
   cu my_cu (inst[31:26], inst[5:0], zero, wmem, wreg, regrt, m2reg,
                        aluc, shift, aluimm, pcsource, jal, sext);

   mux2x32 alu_b (data, immediate, aluimm, alub);
   mux2x32 alu_a (ra, sa, shift, alua);
   mux2x32 result(alu, mem, m2reg, alu_mem);
   mux2x32 link (alu_mem, p4, jal, res);
   mux2x5 reg_wn (inst[15:11], inst[20:16], regrt, reg_dest);
   assign wn = reg_dest | {5{jal}}; // jal: r31 <-- p4;      // 31 or reg_dest
   mux4x32 nextpc(p4, adr, ra, jpc, pcsource, npc);
   regfile rf (inst[25:21], inst[20:16], res, wn, wreg, clock, resetn, ra, data);
   alu al_unit (alua, alub, aluc, alu, zero);
endmodule
